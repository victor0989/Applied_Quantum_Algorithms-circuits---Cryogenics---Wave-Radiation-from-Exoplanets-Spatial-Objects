//Monitoring Temperature And Intensity through IoT with FPGA Device(VHDL) GitHub repository
//Design recipes with FPGA(VHDL) examples 

//Ultrasonic_Sensor.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity Ultrasonic_Sensor is
    port(
       
        pulse_pin in std_logic;
        
        trig_pin: out std_logic;
         rst: in std_logic;

         clk: in std_logic;
         an: out std_logic_vector(2 downto 0);
         sseg: out std_logic_vector (7 downto 0)
       );
end Ultrasonic_Sensor;

arquitectura Behavioral of Ultrasonic_Sensor is

component Range_sensor is
    port(
        fpgaclk, pulse: in std_logic;
        trigger_out: out std_logic;
        meters, decimeters, centimeters: out std_logic_vector(3 downto 0)
);

end component;

compoent display_cts is port
(
  clk: in std_logic;
  Display_reset : in std_logic;
  in2, in1, in0: in std_logic_vector(3) downto 0);
  an: out std_logic_vector(2 downto 0);
  sseg: out std_logic_vector (7 downto 0)
);
end component;

signal Ai: std_logic_vector(3 downto 0);

begin
    range_sens_: Range_sensor port map (clk, puse_pin, trig_pin, Ai, Si, Ci);
display_i; display_ctr port map(clk,rst, Ai,   Bi, Ci,   an,   sseg);

end Behavioral;
